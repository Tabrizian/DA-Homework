package common is
    type gene is (A, T, C, G);
end common;

package body common is
end common;
