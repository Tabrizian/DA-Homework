library ieee;
use ieee.std_logic_1164.all;

package common is
    type array_2d is array (natural) of std_logic_vector(7 downto 0);
end common;
